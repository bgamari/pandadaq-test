`timescale 1ns / 1ps
module pandadaq(
    inout [7:0] ja,
	 output led_red,
	 output led_green,
    inout [7:0] jb,
    output [2:0] ad2_os,
    output ad2_stby,
    output ad2_range,
    output adx_convsta,
    output adx_convstb,
    output adx_reset,
    output adx_sclk,
    output ad2_ncs,
	 input ad2_busy,
    input ad2_douta,
    input ad2_doutb,
    output [2:0] ad1_os,
    output ad1_stby,
    output ad1_range,
    output ad1_ncs,
    input ad1_busy,
    output ad1_douta,
    output ad1_doutb,
    output da_din,
    output da_sclk,
    output da_nldac,
    output da_nsync,
    output fpga_awake,
    output mcspi1_somi,
    input mcspi1_clk,
    input gps_miso,
    output gps_mosi,
    input mcspi1_simo,
    input mcspi1_cs0,
    output gps_on_off,
    output gps_sclk,
    output gps_ncs,
    input gps_1pps,
    inout [7:0] je,
	 input fpga_ocxo,
	 input fpga_clk,
    input fpga_init,
    input mcspi1_cs1,
    inout [15:0] gpmc_ad,
    output gpmc_wait0,
	 inout gpio_54,
    input gpmc_clk,
    input gpmc_nbe0,
    input gpmc_ale,
    input gpmc_ncs0,
    input gpmc_ncs1,
    inout gpio_140,
    input gpmc_noe,
    input gpmc_nwe
    );

blinky blink_green(fpga_clk, led_green);
blinky blink_red(fpga_clk, led_red);

endmodule
